class mult_tlm extends base_tlm#();


endclass : mult_tlm
