`include "base_ifc.sv"
`include "adder_ifc.sv"
`include "mult_ifc.sv"
`include "divider_ifc.sv"
`include "pipeline_ifc.sv"
`include "uart_ifc.sv"

module gpu_tb();

    import gpu_pkg::*;

endmodule
