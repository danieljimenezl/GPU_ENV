interface mult_ifc();

    logic in0_mult [15:0];
    logic in1_mult [15:0];
    logic out_mult [15:0];

endinterface : mult_ifc
