interface adder_ifc();

    logic in0_adder;
    logic in1_adder;
    logic out_adder;

endinterface : adder_ifc    
