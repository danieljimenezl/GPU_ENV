interface adder_ifc();

    base_ifc base();

    logic [15:0] in0_adder;
    logic [15:0] in1_adder;
    logic [15:0] out_adder;

endinterface : adder_ifc    
