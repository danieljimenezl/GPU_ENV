virtual class base_tlm extends uvm_sequence_item;
/*
    `uvm_component_utils_begin(base_tlm)
    `uvm_component_utils_end

    //--------------------------------------------
    // new
    function new (string name);
        super.new(name);
     endfunction : new
*/
endclass : base_tlm
