interface uart_ifc();



endinterface : uart_ifc
