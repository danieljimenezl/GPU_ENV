`include "base_ifc.sv"
`include "adder_ifc.sv"

module gpu_tb();

    import gpu_pkg::*;

endmodule
