class adder_tlm extends base_tlm#();


endclass : adder_tlm
