interface pipeline_ifc();

endinterface : pipeline_ifc    
