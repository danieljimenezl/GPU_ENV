interface pipeline_ifc();

    base_ifc base();

endinterface : pipeline_ifc    
