class divider_tlm extends base_tlm#();


endclass : divider_tlm
