interface divider_ifc();

    base_ifc base();

    logic [15:0] in0_divider;
    logic [15:0] in1_divider;
    logic [15:0] out_divider;

endinterface : divider_ifc
