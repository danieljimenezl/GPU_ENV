package gpu_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    ///////////////////////////////////////////////
    //  G P U - B A S E
    `include "base_seq.sv"
    `include "base_driver.sv"
    `include "base_monitor.sv"
    `include "base_scoreboard.sv"
    //`include "gpu_base/base_agent.sv"

endpackage
