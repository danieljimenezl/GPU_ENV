interface base_ifc();
    logic clk;

endinterface : base_ifc
