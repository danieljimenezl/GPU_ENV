interface divider_ifc();

    logic in0_divider [15:0];
    logic in1_divider [15:0];
    logic out_divider [15:0];

endinterface : divider_ifc
