`include "base_ifc.sv"

module gpu_tb();

    import gpu_pkg::*;

endmodule
