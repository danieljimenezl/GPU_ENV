interface mult_ifc();

    base_ifc base();

    logic [15:0] in0_mult;
    logic [15:0] in1_mult;
    logic [15:0] out_mult;

endinterface : mult_ifc
