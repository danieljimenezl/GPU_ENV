`include "base_ifc.sv"
`include "adder_ifc.sv"
`include "mult_ifc.sv"
`include "divider_ifc.sv"

module gpu_tb();

    import gpu_pkg::*;

endmodule
