interface adder_ifc();

    logic [15:0] in0_adder;
    logic [15:0] in1_adder;
    logic [15:0] out_adder;

endinterface : adder_ifc    
