interface adder_ifc();

    logic in0_adder [15:0];
    logic in1_adder [15:0];
    logic out_adder [15:0];

endinterface : adder_ifc    
